module Execute(
					input wire clock,
					input reg [15:0] r1,
					input reg [15:0] r2,
					input reg [3:0] codop,
					input reg [3:0] imm,
					output reg [15:0] saida_alu
);
endmodule
